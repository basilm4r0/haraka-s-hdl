package harakas_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    typedef uvm_config_db#(virtual harakas_if) harakas_vif_config;

    `include "harakas_message.sv"
    `include "harakas_monitor.sv"
    `include "harakas_sequencer.sv"
    `include "harakas_seqs.sv"
    `include "harakas_driver.sv"
    `include "harakas_agent.sv"
    `include "harakas_scoreboard.sv"
    `include "harakas_env.sv"

endpackage

import uvm_pkg::*;
`include "interface.sv"
`include "sequence_item.sv"
`include "driver.sv"
`include "monitor.sv"
`include "sequencer.sv"
`include "agent.sv"

class haraka_s_sequencer extends uvm_sequencer #(haraka_s_sequence_item);
    
    //1. UVM component
    `uvm_component_utils(haraka_s_sequencer)

    //2. Constructor
    function new(string name = "haraka_s_sequencer", uvm_component parent);
        super.new(name, parent);
    endfunction

    //3. Build Phase
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
    endfunction

endclass: haraka_s_sequencer